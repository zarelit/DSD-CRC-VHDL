-------------------------------------------------------------------------------
--
-- Title       : Configuration preload_conf_crc_control for crc_control
-- Design      : CRCmd
-- Author      : Giuliano
-- Company     : La mia
--
-------------------------------------------------------------------------------
--
-- File        : Z:\DSD\progetto_CRC\CRCmd\src\preload_conf_crc_control.vhd
-- Generated   : 1/10/2013, 2:26 PM
-- From        : no source file
-- By          : Active-HDL Built-in Configuration Generator ver. 1.2s
--
-------------------------------------------------------------------------------
--
-- Description : Automatically generated configuration file for crc_control
--
-------------------------------------------------------------------------------

configuration preload_conf_crc_control of crc_control is
for preload_behave
end for;
end preload_conf_crc_control;
